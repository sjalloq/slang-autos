module top;
    /*AUTOWIRE*/
    // Beginning of automatic wires
    logic old_signal;  // This should be removed
    // End of automatics
    submod u_sub (/*AUTOINST*/);
endmodule
