// Child module with outputs that get consumed by inline wire declaration
module child (
    input  logic clk,
    output logic [3:0] sig_a,
    output logic [3:0] sig_b
);
endmodule
