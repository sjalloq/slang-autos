// Single-bit port module for width adaptation tests
module one_bit(
    input  logic clk,
    input  logic data_in,    // 1-bit input
    output logic data_out    // 1-bit output
);
endmodule
