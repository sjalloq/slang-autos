module top;
    /*AUTOWIRE*/
    /* submod AUTO_TEMPLATE
        data_out => '0
        valid => _
    */
    submod u_sub (/*AUTOINST*/);
endmodule
