module top (
    output logic b
);

    /*AUTOREG*/

    submod u_sub (/*AUTOINST*/);

endmodule