// Test: Packed arrays should preserve structure with resolved-ranges
module top (
    input logic clk
    /*AUTOPORTS*/
);
    /*AUTOLOGIC*/
    child u_child (/*AUTOINST*/);
endmodule
