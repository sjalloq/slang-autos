module top;
    /*AUTOWIRE*/
    /* narrow AUTO_TEMPLATE
        data => shared_bus
    */
    narrow u_narrow (/*AUTOINST*/);
    /* wide AUTO_TEMPLATE
        data => shared_bus
    */
    wide u_wide (/*AUTOINST*/);
endmodule
