module top;
    /*AUTOWIRE*/
    bidir u_bidir (/*AUTOINST*/);
endmodule
