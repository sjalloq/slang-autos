module top;
    // This module does not exist in any library
    nonexistent_module u_missing (/*AUTOINST*/);
endmodule
