module producer (
    input  logic        clk,
    input  logic        rst_n,
    output logic [2:0]  some_sig,    // Drives some_sig
    output logic [7:0]  data_out
);
endmodule
