module debug_module (
    input  logic clk,
    input  logic [31:0] debug_info_l,
    input  logic [31:0] debug_info_h
);
endmodule
