module top
    // Missing semicolon and other syntax errors
    wire clk
    submod u_sub (/*AUTOINST*/)
endmodule
