module submod(
    input logic clk,
    input logic [7:0] data_in,
    output logic [7:0] data_out
);
endmodule
