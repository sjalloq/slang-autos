module submod(
    input wire clk,
    input wire rst_n
);
endmodule
