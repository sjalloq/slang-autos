module top;
    /*AUTOWIRE*/
    submod u_sub (/*AUTOINST*/);
endmodule
