module child3 (
    input  logic clk,
    output logic data_out0,
    output logic data_out1,
    output logic data_out2,
    output logic data_out3
);
endmodule
