module top;
    submod u_sub0 (/*AUTOINST*/);
endmodule
