module top_unsorted (
    input  logic clk,
    input  logic rst_n
    /*AUTOPORTS*/
    output logic valid,
    output logic  [7:0] data_out,
    input logic  [7:0] data_in
);
    /*AUTOWIRE*/

    submod u_sub (/*AUTOINST*/);
endmodule
