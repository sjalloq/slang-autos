module fifo(
    input  wire        clk,
    input  wire        rst_n,
    input  wire [7:0]  din,
    output wire [7:0]  dout,
    output wire        empty,
    output wire        full
);
endmodule
