module submod (
    output logic a
);
endmodule
