// Consumes 8-bit data
module consumer_narrow(
    input  logic       clk,
    input  logic [7:0] data
);
endmodule
