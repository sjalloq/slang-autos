module top;
    logic [7:0] data_out;  // User declared - should be skipped
    /*AUTOWIRE*/
    submod u_sub (/*AUTOINST*/);
endmodule
