module producer (
    input  logic clk,
    output logic [2:0] fifo_level
);
endmodule
