module top;
    /* fifo AUTO_TEMPLATE (
       din  => data_@_in,
       dout => data_@_out,
    ); */
    fifo u_fifo_0 (/*AUTOINST*/);
    fifo u_fifo_1 (/*AUTOINST*/);
endmodule
