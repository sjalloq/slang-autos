module top;
  submod u_sub (/*AUTOINST*/);
endmodule
