module bidir(
    inout logic [7:0] bus
);
endmodule
