// Produces 16-bit data (wider than consumer)
module producer_wide(
    input  logic        clk,
    output logic [15:0] data
);
endmodule
