module child (
    input  logic clk,
    input  logic data_in0,
    input  logic data_in1,
    output logic data_out0,
    output logic data_out1
);
endmodule
