// Child module with multiple inputs
module child (
    input  logic        clk,
    input  logic [3:0]  sig_a,
    input  logic [3:0]  sig_b,
    output logic [7:0]  data_out
);
endmodule
