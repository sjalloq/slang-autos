// Test part select width aggregation
module top_partsel (
    input logic clk
    /*AUTOPORTS*/
);

    /* debug_module AUTO_TEMPLATE
        debug_info_l => cxpl_debug_info[31:0],
        debug_info_h => cxpl_debug_info[63:32],
     */
    debug_module u_debug (/*AUTOINST*/);

endmodule
