// Simple synchronization pulse module for instance array test
module sync_pulse (
    input  logic        clk,
    input  logic        rst_n,
    input  logic [7:0]  data_in,
    output logic [7:0]  data_out,
    output logic        valid
);
    // Synchronization logic
endmodule
