// Consumes 16-bit data (wider than producer)
module consumer_wide(
    input  logic        clk,
    input  logic [15:0] data
);
endmodule
