module submod #(
    parameter WIDTH = 8
)(
    input logic clk,
    input logic [WIDTH-1:0] data_in,
    output logic [WIDTH-1:0] data_out
);
endmodule
