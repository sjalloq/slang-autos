module consumer (
    input  logic        clk,
    input  logic        rst_n,
    input  logic [2:0]  some_sig,    // Receives some_sig
    input  logic [7:0]  data_in
);
endmodule
