// Test: Macro in port widths
`define DATA_WIDTH 8

module top (/*AUTOPORTS*/);
    /*AUTOLOGIC*/
    sub u_sub (/*AUTOINST*/);
endmodule
