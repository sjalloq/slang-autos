// Produces 8-bit data
module producer_narrow(
    input  logic       clk,
    output logic [7:0] data
);
endmodule
