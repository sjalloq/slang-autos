module narrow(
    output logic [7:0] data
);
endmodule
