module child (
    input  logic clk,
    input  logic [2:0] data_in0,
    input  logic [2:0] data_in1,
    input  logic [2:0] data_in2,
    input  logic [2:0] data_in3
);
endmodule
