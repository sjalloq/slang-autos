module top;
    /*AUTOWIRE*/
    /* submod AUTO_TEMPLATE
        data_out => renamed_signal
    */
    submod u_sub (/*AUTOINST*/);
endmodule
