module child (
    input logic a,
    input logic b
);
endmodule
