module child2 (
    input  logic clk,
    input  logic amf_msi_rc_int0_csr_fifo_ovrflw_in,
    input  logic amf_msi_rc_int1_csr_fifo_ovrflw_in,
    input  logic amf_msi_rc_int2_csr_fifo_ovrflw_in,
    input  logic amf_msi_rc_int3_csr_fifo_ovrflw_in
);
endmodule
