module wide(
    output logic [15:0] data
);
endmodule
