// Test: Unpacked arrays should preserve dimensions after signal name
module top (
    input logic clk
    /*AUTOPORTS*/
);
    /*AUTOLOGIC*/
    child u_child (/*AUTOINST*/);
endmodule
